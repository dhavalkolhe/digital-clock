/mnt/c/users/dhava/Desktop/Web-dev/digital-clock